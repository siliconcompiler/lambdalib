module la_pt(a,a);
   inout a;
endmodule // la_pt
