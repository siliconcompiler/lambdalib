
module la_tiehi(z);
  output z;
  sky130_fd_sc_hd__conb_1 _0_ (
    .HI(z)
  );
endmodule
