/*****************************************************************************
 * Function: Padframe Bitfield Definitions
 * Copyright: Lambda Project Authors. ALl rights Reserved.
 * License:  MIT (see LICENSE file in Lambda repository)
 ****************************************************************************/

localparam LA_BIDIR  = 4'h0;
localparam LA_INPUT  = 4'h1;
localparam LA_ANALOG = 4'h2;
localparam LA_XTAL   = 4'h3;
localparam LA_VDDIO  = 4'h8;
localparam LA_VSSIO  = 4'h9;
localparam LA_VDD    = 4'hA;
localparam LA_VSS    = 4'hB;
localparam LA_VDDA   = 4'hC;
localparam LA_VSSA   = 4'hD;
localparam LA_POC    = 4'hE;
localparam LA_CUT    = 4'hF;
