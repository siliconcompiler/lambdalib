/*****************************************************************************
 * Function: IO bidirectional buffer
 * Copyright: Lambda Project Authors. ALl rights Reserved.
 * License:  MIT (see LICENSE file in Lambda repository)
 *
 * Docs:
 * This is a generic cell that defines the standard interface of the lambda
 * bidrectional buffer cell. It is only suitable for FPGA synthesis.
 *
 * ASIC specific libraries will need to use the TYPE field to select an
 * appropriate hardcoded physical cell based on the the process constraints
 * and library composition. For example, modern nodes will usually have
 * different IP cells for the placing cells vvertically or horizontally.
 *
 ****************************************************************************/
module la_iobidir
  #(
    parameter TYPE = "DEFAULT" // cell type
    )
   (// io pad signals
    inout 	 pad, // bidirectional pad signal
    inout 	 vdd, // core supply
    inout 	 vss, // core ground
    inout 	 vddio, // io supply
    inout 	 vssio, // io ground
    // core facing signals
    input 	 a, // input from core
    output 	 z, // output to core
    input 	 ie, // input enable, 1 = active
    input 	 oe, // output enable, 1 = active
    input 	 pe, // weak pull enable, 1 = active
    input 	 ps,// pull select, 1 = pull-up, 0 = pull-down
    input 	 sr, // slewrate enable 1 = fast, 0 = slow
    input [2:0]  ds, // drive strength, 3'b0 = weakest
    input 	 st, // schmitt trigger, 1 = enable
    inout [7:0]  ioring, // generic io-ring interface
    input [31:0] cfg // generic config interface
    );

   // to core
   assign z   = ie ? pad : 1'b0;

   // to pad (verilator only)
   assign pad = oe         ? a    :
		(pe & ps)  ? 1'b1 :
		(pe & !ps) ? 1'b0 :
                             1'bz;

endmodule
