
module la_delay(a, z);
  input a;
  output z;
  assign z = a;
endmodule
