/*****************************************************************************
 * Function: Padring Generator Enumeration
 * Copyright: Lambda Project Authors. All rights Reserved.
 * License:  MIT (see LICENSE file in Lambda repository)
 ****************************************************************************/

// NULL (place holder)
localparam [7:0] NULL      = 8'h00;

// io cells
localparam [7:0] LA_BIDIR  = 8'h01;
localparam [7:0] LA_INPUT  = 8'h02;
localparam [7:0] LA_OUTPUT = 8'h03;
localparam [7:0] LA_ANALOG = 8'h04;
localparam [7:0] LA_XTAL   = 8'h05;
localparam [7:0] LA_RXDIFF = 8'h06;
localparam [7:0] LA_TXDIFF = 8'h07;

// supply cells
localparam [7:0] LA_VDDIO  = 8'h10;
localparam [7:0] LA_VSSIO  = 8'h11;
localparam [7:0] LA_VDD    = 8'h12;
localparam [7:0] LA_VSS    = 8'h13;
localparam [7:0] LA_VDDA   = 8'h14;
localparam [7:0] LA_VSSA   = 8'h15;
localparam [7:0] LA_POC    = 8'h16;
localparam [7:0] LA_CUT    = 8'h17;
localparam [7:0] LA_CLAMP  = 8'h18;

// simple pin enumeration
localparam [7:0] PIN0  = 8'd00;
localparam [7:0] PIN1  = 8'd01;
localparam [7:0] PIN2  = 8'd02;
localparam [7:0] PIN3  = 8'd03;
localparam [7:0] PIN4  = 8'd04;
localparam [7:0] PIN5  = 8'd05;
localparam [7:0] PIN6  = 8'd06;
localparam [7:0] PIN7  = 8'd07;
localparam [7:0] PIN8  = 8'd08;
localparam [7:0] PIN9  = 8'd09;
localparam [7:0] PIN10 = 8'd10;
localparam [7:0] PIN11 = 8'd11;
localparam [7:0] PIN12 = 8'd12;
localparam [7:0] PIN13 = 8'd13;
localparam [7:0] PIN14 = 8'd14;
localparam [7:0] PIN15 = 8'd15;

localparam [7:0] PIN16 = 8'd16;
localparam [7:0] PIN17 = 8'd17;
localparam [7:0] PIN18 = 8'd18;
localparam [7:0] PIN19 = 8'd19;
localparam [7:0] PIN20 = 8'd20;
localparam [7:0] PIN21 = 8'd21;
localparam [7:0] PIN22 = 8'd22;
localparam [7:0] PIN23 = 8'd23;
localparam [7:0] PIN24 = 8'd24;
localparam [7:0] PIN25 = 8'd25;
localparam [7:0] PIN26 = 8'd26;
localparam [7:0] PIN27 = 8'd27;
localparam [7:0] PIN28 = 8'd28;
localparam [7:0] PIN29 = 8'd29;
localparam [7:0] PIN30 = 8'd30;
localparam [7:0] PIN31 = 8'd31;

localparam [7:0] PIN32 = 8'd32;
localparam [7:0] PIN33 = 8'd33;
localparam [7:0] PIN34 = 8'd34;
localparam [7:0] PIN35 = 8'd35;
localparam [7:0] PIN36 = 8'd36;
localparam [7:0] PIN37 = 8'd37;
localparam [7:0] PIN38 = 8'd38;
localparam [7:0] PIN39 = 8'd39;
localparam [7:0] PIN40 = 8'd40;
localparam [7:0] PIN41 = 8'd41;
localparam [7:0] PIN42 = 8'd42;
localparam [7:0] PIN43 = 8'd43;
localparam [7:0] PIN44 = 8'd44;
localparam [7:0] PIN45 = 8'd45;
localparam [7:0] PIN46 = 8'd46;
localparam [7:0] PIN47 = 8'd47;

localparam [7:0] PIN48 = 8'd48;
localparam [7:0] PIN49 = 8'd49;
localparam [7:0] PIN50 = 8'd50;
localparam [7:0] PIN51 = 8'd51;
localparam [7:0] PIN52 = 8'd52;
localparam [7:0] PIN53 = 8'd53;
localparam [7:0] PIN54 = 8'd54;
localparam [7:0] PIN55 = 8'd55;
localparam [7:0] PIN56 = 8'd56;
localparam [7:0] PIN57 = 8'd57;
localparam [7:0] PIN58 = 8'd58;
localparam [7:0] PIN59 = 8'd59;
localparam [7:0] PIN60 = 8'd60;
localparam [7:0] PIN61 = 8'd61;
localparam [7:0] PIN62 = 8'd62;
localparam [7:0] PIN63 = 8'd63;
