
module la_clkbuf(a, z);
  input a;
  output z;
  assign z = a;
endmodule
