
module la_tbuf(a, oe, z);
  input a;
  input oe;
  output z;
  assign z = a;
endmodule
