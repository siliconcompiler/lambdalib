/*****************************************************************************
 * Function: 4-Bit Look-Up-Table
 * Copyright: Lambda Project Authors. All rights Reserved.
 * License:  MIT (see LICENSE file in Lambda repository)
 ****************************************************************************/

module la_lut4
  #(parameter TYPE  = "DEFAULT", //  implementation selector
    )
   (input        i0,
    input        i1,
    input        i2,
    input        i3,
    input [15:0] lut,
    output       out
    );

   // 16:8

   // 8:4

   // 4:2

   // 2:1


endmodule
