
module la_tielo(z);
  output z;
  sky130_fd_sc_hd__conb_1 _0_ (
    .LO(z)
  );
endmodule
