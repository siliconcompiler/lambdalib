//#############################################################################
//# Function: And-Or-Inverter (aoi211) Gate                                   #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

module la_aoi211 #(
    parameter PROP = "DEFAULT"
) (
    input  a0,
    input  a1,
    input  b0,
    input  c0,
    output z
);

    assign z = ~((a0 & a1) | b0 | c0);

endmodule
