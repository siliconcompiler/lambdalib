
module la_buf(a, z);
  input a;
  output z;
  assign z = a;
endmodule
