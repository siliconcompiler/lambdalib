//#############################################################################
//# Function: Positive edge-triggered static D-type flop-flop with scan input #
//#                                                                           #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

module la_sdffq #(parameter PROP = "DEFAULT")   (
    input      d,
    input      si,
    input      se,
    input      clk,
    output reg q
    );

   always @ (posedge clk)
       q <= se ? si : d;

endmodule
