/*****************************************************************************
 * Function: Padframe Bitfield Definitions
 * Copyright: Lambda Project Authors. All rights Reserved.
 * License:  MIT (see LICENSE file in Lambda repository)
 ****************************************************************************/

localparam LA_BIDIR = 8'h00;
localparam LA_INPUT = 8'h01;
localparam LA_ANALOG = 8'h02;
localparam LA_XTAL = 8'h03;
localparam LA_VDDIO = 8'h08;
localparam LA_VSSIO = 8'h09;
localparam LA_VDD = 8'h0A;
localparam LA_VSS = 8'h0B;
localparam LA_VDDA = 8'h0C;
localparam LA_VSSA = 8'h0D;
localparam LA_POC = 8'h0E;
localparam LA_CUT = 8'h0F;
localparam LA_DUMMY = 8'h07;
