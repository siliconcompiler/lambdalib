//#############################################################################
//# Function: 2-Input AND Gate                                                #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

module la_and2 #(parameter PROP = "DEFAULT")  (
   input  a,
   input  b,
   output z
   );

   assign z = a & b;

endmodule
