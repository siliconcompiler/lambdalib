//#############################################################################
//# Function: Tie Low Cell                                                    #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

module la_tielo #(
    parameter PROP = "DEFAULT"
) (
    output z
);

    assign z = 1'b0;

endmodule
