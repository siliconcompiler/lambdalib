module sram();

   // TODO: put in la_spram

endmodule
