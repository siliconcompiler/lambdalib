//#############################################################################
//# Function: Tie High Cell                                                   #
//# Copyright: Lambda Project Authors. All rights Reserved.                   #
//# License:  MIT (see LICENSE file in Lambda repository)                     #
//#############################################################################

module la_tiehi #(
    parameter PROP = "DEFAULT"
) (
    output z
);

    assign z = 1'b1;

endmodule
